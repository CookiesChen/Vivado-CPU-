`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/05/24 01:48:24
// Design Name: 
// Module Name: Choose_reg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Choose_reg(
    input ALUSrcA,
    input ALUSrcB,
    input [31:0] ReadData1,
    input [4:0] sa,
    input [31:0] ReadData2,
    input [31:0] exten,
    output [31:0] rega,
    output [31:0] regb
    );
    
    
    
    
endmodule
